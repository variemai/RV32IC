`include "PipelineRegs.v"
module decoder(
    input clk,
    input reset,
    input PipelineRegs::ID_STATE,
    output PipelineRegs::EX_STATE
    );

endmodule
