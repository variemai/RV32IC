program RegisterFile_test(
	input clk,
	output logic we,
	output logic [4:0] read_addr0,
	output logic [4:0] read_addr1,
	output logic [4:0] write_addr,
	output logic [31:0] din,
	input logic [31:0] dout0,
	input logic [31:0] dout1
);
	logic [4:0] ra1 = 5'b0;
	logic [4:0] ra2 = 5'b1;
	logic [31:0] write_data = 8'h0000ffff;
	integer i;
	initial begin
		for(i=0; i<30; i++) begin
			read();
			ra1 = ra1 + 1;
			ra2 = ra2 + 1;
		end
		ra1 = 5'b0;
		ra2 = 5'b1;
		for(i=0; i<30; i++) begin
			$write("ReadWrite\n");
			readwrite();
			ra1 = ra1 + 1;
			ra2 = ra2 + 1;
			write_data = write_data + 1;
		end
		ra1 = 5'b0;
		ra2 = 5'b1;
		for(i=0; i<30; i++) begin
			read();
			ra1 = ra1 + 1;
			ra2 = ra2 + 1;
		end
	end

	task read();
		$write("READ ADDR: %d %d\n",ra1,ra2);
		@(posedge clk) begin
			read_addr0 <= ra1;
			read_addr1 <= ra2;
		end
		@(posedge clk) begin
			$write("DOUT0: %x\n",dout0);
			$write("DOUT1: %x\n",dout1);
		end
	endtask

	task write();
		$write("WRITE ADDR: %d\n",ra1);
		@(posedge clk) begin
			write_addr <= ra1;
			din <= ra2;
			we <= 1;
		end
		@(posedge clk) begin
			we <= 0;
		end
	endtask

	task readwrite();
		@(posedge clk) begin
			write_addr <= ra1;
			we <= 1;
			din <= write_data;
			read_addr0 <= ra1;
			read_addr1 <= ra2;
		end
		@(posedge clk) begin
			we <= 0;
			assert(dout0 == write_data) else 
			$write("DOUT0: %x\n",dout0);
			//$write("DOUT1: %x\n",dout1);
		end
	endtask

endprogram
