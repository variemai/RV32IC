/*****************************************************************************
 * The RV32I Base Instruction Set opcodes as is defined in                   *
 * Volume I: RISC-V User-Level ISA V2.2                                      *
 * Authors: Vardas Ioannis                                                   *
 * created for the purposes of CS-523 RISC-V 32 bit implementation project   *
 * Computer Science Department University of Crete 27/03/2018                *
 *****************************************************************************/

package BIS;
    `define LUI 32'b?????????????????????????0110111
    `define AUIPC 32'b?????????????????????????0010111
    `define JAL 32'b?????????????????????????1101111
    `define JALR 32'b?????????????????000?????1100111
    `define BEQ 32'b????????????????000??????1100011
    `define BNE 32'b????????????????001??????1100011
    `define BLT 32'b????????????????100??????1100011
    `define BGE 32'b????????????????101??????1100011
    `define BLTU 32'b????????????????110??????1100011
    `define BGEU 32'b????????????????111??????1100011
    `define LB 32'b?????????????????000?????0000011
    `define LH 32'b?????????????????001?????0000011
    `define LW 32'b?????????????????010?????0000011
    `define LBU 32'b?????????????????100?????0000011
    `define LHU 32'b?????????????????101?????0000011
endpackage
