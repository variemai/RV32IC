`ifndef _INSTRUCTIONS_SV_
`define _INSTRUCTIONS_SV_

package Instructions;
	`define ILL 16'b0000000000000000
	`define C_ADDI4SPN 16'b000???????????00 	//RES, nzuimm=0
	`define C_LW 16'b010???????????00
	`define C_SW 16'b110???????????00
	`define C_NOP 16'b0000000000000001
	`define C_ADDI 16'b000???????????01 	//HINT, nzimm=0
	`define C_JAL 16'b001???????????01
	`define C_LI 16'b010???????????01 	//HINT, rd=0
	`define C_ADDI16SP 16'b011?00010?????01 	//RES, nzimm=0
	`define C_LUI 16'b011???????????01 	//RES, nzimm=0; HINT, rd=0
	`define C_SRLI 16'b100?00????????01 	//NSE, nzuimm[5]=1
	`define C_SRLI64 16'b100000???0000001 	//ASK FOR DETAILS!!!, HINT 
	`define C_SRAI 16'b100?01????????01	//NSE, nzuimm[5]=1
	`define C_SRAI64 16'b100001???0000001	//ASK FOR DETAILS!!!, HINT
	`define C_ANDI 16'b100?10????????01
	`define C_SUB 16'b100011???00???01
	`define C_XOR 16'b100011???01???01
	`define C_OR 16'b100011???10???01
	`define C_AND 16'b100011???11???01
	`define C_J 16'b101???????????01
	`define C_BEQZ 16'b110???????????01
	`define C_BNEZ 16'b111???????????01
	`define C_SLLI 16'b000???????????10	// HINT, rd=0; NSE, nzuimm[5]=1,
	`define C_SLLI64 16'b0000?????0000010	//HINT
	`define C_LWSP 16'b010???????????10	//RES, rd=0
	`define C_JR 16'b1000?????0000010	//RES, rs1=0
	`define C_MV 16'b1000??????????10	//HINT, rd=0
	`define C_EBREAK 16'b1001000000000010
	`define C_JALR 16'b1001?????0000010
	`define C_ADD 16'b1001??????????10	//HINT, rd=0
	`define C_SWSP 16'b110???????????10

//custom-0 instruction set --> instruction[6:0] = 7'b0001011
//custom-1 instruction set --> instruction[6:0] = 7'b0101011

//`define C.FLD		16'b001???????????00	//RV32DC-only
//`define C.FLW		16'b011???????????00	//RV32FC-only
//`define 			16'b100-----------00	//Reserved
//`define C.FSD		16'b101???????????00	//RV32DC-only
//`define C.FSW		16'b111???????????00	//RV32FC-only
//`define 			16'b100111---10---01	//Reserved
//`define			16'b100111---11---01	//Reserved
//`define C.FLDSP	16'b001???????????10	//RV32DC-only
//`define C.FLWSP	16'b011???????????10	//RV32FC-only
//`define C.FSDSP	16'b101???????????10	//RV32DC-only
//`define C.FSWSP	16'b111???????????10	//RV32FC-only
endpackage
`endif
